module sine_synth (
    input clk,  // clock, 50 Mhz
    input [9:0]FTV,  // frequency tuning value
    input rst,  // reset
    output reg [11:0]dataOut  
  );


  parameter tableSize = 10;
  parameter countSize = 17;
  wire [tableSize-1:0]prioBits;
  reg [countSize-1:0]counter; 
  
  //store half the table size
  wire [11:0] sineval [511:0];
  /* Sequential Logic */
  always @(posedge clk) begin
    if (rst) begin
      counter <= 0;
    end 
    else begin
      counter <= counter + FTV;
    end
    if(prioBits < 512)
      dataOut <= sineval[prioBits];
    else
      dataOut <= 4095-sineval[prioBits-512];
  end
  
  //we have our table size as 10 bits, but in reality,
  //we only store half of the table
  /* Combinational Logic */
  assign prioBits = counter[countSize-1:(countSize-1)-(tableSize-1)];
  
  assign sineval[0] = 2048;
  assign sineval[1] = 2060;
  assign sineval[2] = 2072;
  assign sineval[3] = 2085;
  assign sineval[4] = 2097;
  assign sineval[5] = 2110;
  assign sineval[6] = 2122;
  assign sineval[7] = 2135;
  assign sineval[8] = 2147;
  assign sineval[9] = 2160;
  assign sineval[10] = 2173;
  assign sineval[11] = 2185;
  assign sineval[12] = 2198;
  assign sineval[13] = 2210;
  assign sineval[14] = 2223;
  assign sineval[15] = 2235;
  assign sineval[16] = 2248;
  assign sineval[17] = 2260;
  assign sineval[18] = 2273;
  assign sineval[19] = 2285;
  assign sineval[20] = 2298;
  assign sineval[21] = 2310;
  assign sineval[22] = 2322;
  assign sineval[23] = 2335;
  assign sineval[24] = 2347;
  assign sineval[25] = 2360;
  assign sineval[26] = 2372;
  assign sineval[27] = 2385;
  assign sineval[28] = 2397;
  assign sineval[29] = 2409;
  assign sineval[30] = 2422;
  assign sineval[31] = 2434;
  assign sineval[32] = 2446;
  assign sineval[33] = 2459;
  assign sineval[34] = 2471;
  assign sineval[35] = 2483;
  assign sineval[36] = 2496;
  assign sineval[37] = 2508;
  assign sineval[38] = 2520;
  assign sineval[39] = 2532;
  assign sineval[40] = 2544;
  assign sineval[41] = 2557;
  assign sineval[42] = 2569;
  assign sineval[43] = 2581;
  assign sineval[44] = 2593;
  assign sineval[45] = 2605;
  assign sineval[46] = 2617;
  assign sineval[47] = 2629;
  assign sineval[48] = 2641;
  assign sineval[49] = 2653;
  assign sineval[50] = 2665;
  assign sineval[51] = 2677;
  assign sineval[52] = 2689;
  assign sineval[53] = 2701;
  assign sineval[54] = 2713;
  assign sineval[55] = 2725;
  assign sineval[56] = 2737;
  assign sineval[57] = 2748;
  assign sineval[58] = 2760;
  assign sineval[59] = 2772;
  assign sineval[60] = 2784;
  assign sineval[61] = 2795;
  assign sineval[62] = 2807;
  assign sineval[63] = 2819;
  assign sineval[64] = 2830;
  assign sineval[65] = 2842;
  assign sineval[66] = 2854;
  assign sineval[67] = 2865;
  assign sineval[68] = 2877;
  assign sineval[69] = 2888;
  assign sineval[70] = 2899;
  assign sineval[71] = 2911;
  assign sineval[72] = 2922;
  assign sineval[73] = 2934;
  assign sineval[74] = 2945;
  assign sineval[75] = 2956;
  assign sineval[76] = 2967;
  assign sineval[77] = 2979;
  assign sineval[78] = 2990;
  assign sineval[79] = 3001;
  assign sineval[80] = 3012;
  assign sineval[81] = 3023;
  assign sineval[82] = 3034;
  assign sineval[83] = 3045;
  assign sineval[84] = 3056;
  assign sineval[85] = 3067;
  assign sineval[86] = 3078;
  assign sineval[87] = 3089;
  assign sineval[88] = 3099;
  assign sineval[89] = 3110;
  assign sineval[90] = 3121;
  assign sineval[91] = 3132;
  assign sineval[92] = 3142;
  assign sineval[93] = 3153;
  assign sineval[94] = 3163;
  assign sineval[95] = 3174;
  assign sineval[96] = 3184;
  assign sineval[97] = 3195;
  assign sineval[98] = 3205;
  assign sineval[99] = 3215;
  assign sineval[100] = 3226;
  assign sineval[101] = 3236;
  assign sineval[102] = 3246;
  assign sineval[103] = 3256;
  assign sineval[104] = 3266;
  assign sineval[105] = 3276;
  assign sineval[106] = 3286;
  assign sineval[107] = 3296;
  assign sineval[108] = 3306;
  assign sineval[109] = 3316;
  assign sineval[110] = 3326;
  assign sineval[111] = 3336;
  assign sineval[112] = 3346;
  assign sineval[113] = 3355;
  assign sineval[114] = 3365;
  assign sineval[115] = 3375;
  assign sineval[116] = 3384;
  assign sineval[117] = 3394;
  assign sineval[118] = 3403;
  assign sineval[119] = 3412;
  assign sineval[120] = 3422;
  assign sineval[121] = 3431;
  assign sineval[122] = 3440;
  assign sineval[123] = 3449;
  assign sineval[124] = 3458;
  assign sineval[125] = 3468;
  assign sineval[126] = 3477;
  assign sineval[127] = 3486;
  assign sineval[128] = 3494;
  assign sineval[129] = 3503;
  assign sineval[130] = 3512;
  assign sineval[131] = 3521;
  assign sineval[132] = 3530;
  assign sineval[133] = 3538;
  assign sineval[134] = 3547;
  assign sineval[135] = 3555;
  assign sineval[136] = 3564;
  assign sineval[137] = 3572;
  assign sineval[138] = 3580;
  assign sineval[139] = 3589;
  assign sineval[140] = 3597;
  assign sineval[141] = 3605;
  assign sineval[142] = 3613;
  assign sineval[143] = 3621;
  assign sineval[144] = 3629;
  assign sineval[145] = 3637;
  assign sineval[146] = 3645;
  assign sineval[147] = 3653;
  assign sineval[148] = 3661;
  assign sineval[149] = 3668;
  assign sineval[150] = 3676;
  assign sineval[151] = 3684;
  assign sineval[152] = 3691;
  assign sineval[153] = 3699;
  assign sineval[154] = 3706;
  assign sineval[155] = 3713;
  assign sineval[156] = 3721;
  assign sineval[157] = 3728;
  assign sineval[158] = 3735;
  assign sineval[159] = 3742;
  assign sineval[160] = 3749;
  assign sineval[161] = 3756;
  assign sineval[162] = 3763;
  assign sineval[163] = 3770;
  assign sineval[164] = 3776;
  assign sineval[165] = 3783;
  assign sineval[166] = 3790;
  assign sineval[167] = 3796;
  assign sineval[168] = 3803;
  assign sineval[169] = 3809;
  assign sineval[170] = 3816;
  assign sineval[171] = 3822;
  assign sineval[172] = 3828;
  assign sineval[173] = 3834;
  assign sineval[174] = 3840;
  assign sineval[175] = 3846;
  assign sineval[176] = 3852;
  assign sineval[177] = 3858;
  assign sineval[178] = 3864;
  assign sineval[179] = 3870;
  assign sineval[180] = 3875;
  assign sineval[181] = 3881;
  assign sineval[182] = 3887;
  assign sineval[183] = 3892;
  assign sineval[184] = 3897;
  assign sineval[185] = 3903;
  assign sineval[186] = 3908;
  assign sineval[187] = 3913;
  assign sineval[188] = 3918;
  assign sineval[189] = 3923;
  assign sineval[190] = 3928;
  assign sineval[191] = 3933;
  assign sineval[192] = 3938;
  assign sineval[193] = 3943;
  assign sineval[194] = 3948;
  assign sineval[195] = 3952;
  assign sineval[196] = 3957;
  assign sineval[197] = 3961;
  assign sineval[198] = 3966;
  assign sineval[199] = 3970;
  assign sineval[200] = 3974;
  assign sineval[201] = 3979;
  assign sineval[202] = 3983;
  assign sineval[203] = 3987;
  assign sineval[204] = 3991;
  assign sineval[205] = 3995;
  assign sineval[206] = 3998;
  assign sineval[207] = 4002;
  assign sineval[208] = 4006;
  assign sineval[209] = 4009;
  assign sineval[210] = 4013;
  assign sineval[211] = 4016;
  assign sineval[212] = 4020;
  assign sineval[213] = 4023;
  assign sineval[214] = 4026;
  assign sineval[215] = 4030;
  assign sineval[216] = 4033;
  assign sineval[217] = 4036;
  assign sineval[218] = 4039;
  assign sineval[219] = 4041;
  assign sineval[220] = 4044;
  assign sineval[221] = 4047;
  assign sineval[222] = 4050;
  assign sineval[223] = 4052;
  assign sineval[224] = 4055;
  assign sineval[225] = 4057;
  assign sineval[226] = 4059;
  assign sineval[227] = 4062;
  assign sineval[228] = 4064;
  assign sineval[229] = 4066;
  assign sineval[230] = 4068;
  assign sineval[231] = 4070;
  assign sineval[232] = 4072;
  assign sineval[233] = 4074;
  assign sineval[234] = 4075;
  assign sineval[235] = 4077;
  assign sineval[236] = 4079;
  assign sineval[237] = 4080;
  assign sineval[238] = 4082;
  assign sineval[239] = 4083;
  assign sineval[240] = 4084;
  assign sineval[241] = 4085;
  assign sineval[242] = 4086;
  assign sineval[243] = 4087;
  assign sineval[244] = 4088;
  assign sineval[245] = 4089;
  assign sineval[246] = 4090;
  assign sineval[247] = 4091;
  assign sineval[248] = 4092;
  assign sineval[249] = 4092;
  assign sineval[250] = 4093;
  assign sineval[251] = 4093;
  assign sineval[252] = 4093;
  assign sineval[253] = 4094;
  assign sineval[254] = 4094;
  assign sineval[255] = 4094;
  assign sineval[256] = 4094;
  assign sineval[257] = 4094;
  assign sineval[258] = 4094;
  assign sineval[259] = 4094;
  assign sineval[260] = 4093;
  assign sineval[261] = 4093;
  assign sineval[262] = 4093;
  assign sineval[263] = 4092;
  assign sineval[264] = 4092;
  assign sineval[265] = 4091;
  assign sineval[266] = 4090;
  assign sineval[267] = 4089;
  assign sineval[268] = 4088;
  assign sineval[269] = 4087;
  assign sineval[270] = 4086;
  assign sineval[271] = 4085;
  assign sineval[272] = 4084;
  assign sineval[273] = 4083;
  assign sineval[274] = 4082;
  assign sineval[275] = 4080;
  assign sineval[276] = 4079;
  assign sineval[277] = 4077;
  assign sineval[278] = 4075;
  assign sineval[279] = 4074;
  assign sineval[280] = 4072;
  assign sineval[281] = 4070;
  assign sineval[282] = 4068;
  assign sineval[283] = 4066;
  assign sineval[284] = 4064;
  assign sineval[285] = 4062;
  assign sineval[286] = 4059;
  assign sineval[287] = 4057;
  assign sineval[288] = 4055;
  assign sineval[289] = 4052;
  assign sineval[290] = 4050;
  assign sineval[291] = 4047;
  assign sineval[292] = 4044;
  assign sineval[293] = 4041;
  assign sineval[294] = 4039;
  assign sineval[295] = 4036;
  assign sineval[296] = 4033;
  assign sineval[297] = 4030;
  assign sineval[298] = 4026;
  assign sineval[299] = 4023;
  assign sineval[300] = 4020;
  assign sineval[301] = 4016;
  assign sineval[302] = 4013;
  assign sineval[303] = 4009;
  assign sineval[304] = 4006;
  assign sineval[305] = 4002;
  assign sineval[306] = 3998;
  assign sineval[307] = 3995;
  assign sineval[308] = 3991;
  assign sineval[309] = 3987;
  assign sineval[310] = 3983;
  assign sineval[311] = 3979;
  assign sineval[312] = 3974;
  assign sineval[313] = 3970;
  assign sineval[314] = 3966;
  assign sineval[315] = 3961;
  assign sineval[316] = 3957;
  assign sineval[317] = 3952;
  assign sineval[318] = 3948;
  assign sineval[319] = 3943;
  assign sineval[320] = 3938;
  assign sineval[321] = 3933;
  assign sineval[322] = 3928;
  assign sineval[323] = 3923;
  assign sineval[324] = 3918;
  assign sineval[325] = 3913;
  assign sineval[326] = 3908;
  assign sineval[327] = 3903;
  assign sineval[328] = 3897;
  assign sineval[329] = 3892;
  assign sineval[330] = 3887;
  assign sineval[331] = 3881;
  assign sineval[332] = 3875;
  assign sineval[333] = 3870;
  assign sineval[334] = 3864;
  assign sineval[335] = 3858;
  assign sineval[336] = 3852;
  assign sineval[337] = 3846;
  assign sineval[338] = 3840;
  assign sineval[339] = 3834;
  assign sineval[340] = 3828;
  assign sineval[341] = 3822;
  assign sineval[342] = 3816;
  assign sineval[343] = 3809;
  assign sineval[344] = 3803;
  assign sineval[345] = 3796;
  assign sineval[346] = 3790;
  assign sineval[347] = 3783;
  assign sineval[348] = 3776;
  assign sineval[349] = 3770;
  assign sineval[350] = 3763;
  assign sineval[351] = 3756;
  assign sineval[352] = 3749;
  assign sineval[353] = 3742;
  assign sineval[354] = 3735;
  assign sineval[355] = 3728;
  assign sineval[356] = 3721;
  assign sineval[357] = 3713;
  assign sineval[358] = 3706;
  assign sineval[359] = 3699;
  assign sineval[360] = 3691;
  assign sineval[361] = 3684;
  assign sineval[362] = 3676;
  assign sineval[363] = 3668;
  assign sineval[364] = 3661;
  assign sineval[365] = 3653;
  assign sineval[366] = 3645;
  assign sineval[367] = 3637;
  assign sineval[368] = 3629;
  assign sineval[369] = 3621;
  assign sineval[370] = 3613;
  assign sineval[371] = 3605;
  assign sineval[372] = 3597;
  assign sineval[373] = 3589;
  assign sineval[374] = 3580;
  assign sineval[375] = 3572;
  assign sineval[376] = 3564;
  assign sineval[377] = 3555;
  assign sineval[378] = 3547;
  assign sineval[379] = 3538;
  assign sineval[380] = 3530;
  assign sineval[381] = 3521;
  assign sineval[382] = 3512;
  assign sineval[383] = 3503;
  assign sineval[384] = 3494;
  assign sineval[385] = 3486;
  assign sineval[386] = 3477;
  assign sineval[387] = 3468;
  assign sineval[388] = 3458;
  assign sineval[389] = 3449;
  assign sineval[390] = 3440;
  assign sineval[391] = 3431;
  assign sineval[392] = 3422;
  assign sineval[393] = 3412;
  assign sineval[394] = 3403;
  assign sineval[395] = 3394;
  assign sineval[396] = 3384;
  assign sineval[397] = 3375;
  assign sineval[398] = 3365;
  assign sineval[399] = 3355;
  assign sineval[400] = 3346;
  assign sineval[401] = 3336;
  assign sineval[402] = 3326;
  assign sineval[403] = 3316;
  assign sineval[404] = 3306;
  assign sineval[405] = 3296;
  assign sineval[406] = 3286;
  assign sineval[407] = 3276;
  assign sineval[408] = 3266;
  assign sineval[409] = 3256;
  assign sineval[410] = 3246;
  assign sineval[411] = 3236;
  assign sineval[412] = 3226;
  assign sineval[413] = 3215;
  assign sineval[414] = 3205;
  assign sineval[415] = 3195;
  assign sineval[416] = 3184;
  assign sineval[417] = 3174;
  assign sineval[418] = 3163;
  assign sineval[419] = 3153;
  assign sineval[420] = 3142;
  assign sineval[421] = 3132;
  assign sineval[422] = 3121;
  assign sineval[423] = 3110;
  assign sineval[424] = 3099;
  assign sineval[425] = 3089;
  assign sineval[426] = 3078;
  assign sineval[427] = 3067;
  assign sineval[428] = 3056;
  assign sineval[429] = 3045;
  assign sineval[430] = 3034;
  assign sineval[431] = 3023;
  assign sineval[432] = 3012;
  assign sineval[433] = 3001;
  assign sineval[434] = 2990;
  assign sineval[435] = 2979;
  assign sineval[436] = 2967;
  assign sineval[437] = 2956;
  assign sineval[438] = 2945;
  assign sineval[439] = 2934;
  assign sineval[440] = 2922;
  assign sineval[441] = 2911;
  assign sineval[442] = 2899;
  assign sineval[443] = 2888;
  assign sineval[444] = 2877;
  assign sineval[445] = 2865;
  assign sineval[446] = 2854;
  assign sineval[447] = 2842;
  assign sineval[448] = 2830;
  assign sineval[449] = 2819;
  assign sineval[450] = 2807;
  assign sineval[451] = 2795;
  assign sineval[452] = 2784;
  assign sineval[453] = 2772;
  assign sineval[454] = 2760;
  assign sineval[455] = 2748;
  assign sineval[456] = 2737;
  assign sineval[457] = 2725;
  assign sineval[458] = 2713;
  assign sineval[459] = 2701;
  assign sineval[460] = 2689;
  assign sineval[461] = 2677;
  assign sineval[462] = 2665;
  assign sineval[463] = 2653;
  assign sineval[464] = 2641;
  assign sineval[465] = 2629;
  assign sineval[466] = 2617;
  assign sineval[467] = 2605;
  assign sineval[468] = 2593;
  assign sineval[469] = 2581;
  assign sineval[470] = 2569;
  assign sineval[471] = 2557;
  assign sineval[472] = 2544;
  assign sineval[473] = 2532;
  assign sineval[474] = 2520;
  assign sineval[475] = 2508;
  assign sineval[476] = 2496;
  assign sineval[477] = 2483;
  assign sineval[478] = 2471;
  assign sineval[479] = 2459;
  assign sineval[480] = 2446;
  assign sineval[481] = 2434;
  assign sineval[482] = 2422;
  assign sineval[483] = 2409;
  assign sineval[484] = 2397;
  assign sineval[485] = 2385;
  assign sineval[486] = 2372;
  assign sineval[487] = 2360;
  assign sineval[488] = 2347;
  assign sineval[489] = 2335;
  assign sineval[490] = 2322;
  assign sineval[491] = 2310;
  assign sineval[492] = 2298;
  assign sineval[493] = 2285;
  assign sineval[494] = 2273;
  assign sineval[495] = 2260;
  assign sineval[496] = 2248;
  assign sineval[497] = 2235;
  assign sineval[498] = 2223;
  assign sineval[499] = 2210;
  assign sineval[500] = 2198;
  assign sineval[501] = 2185;
  assign sineval[502] = 2173;
  assign sineval[503] = 2160;
  assign sineval[504] = 2147;
  assign sineval[505] = 2135;
  assign sineval[506] = 2122;
  assign sineval[507] = 2110;
  assign sineval[508] = 2097;
  assign sineval[509] = 2085;
  assign sineval[510] = 2072;
  assign sineval[511] = 2060;
  
  /*
  always @* begin
   case(prioBits)
			 0 : dataOut   <= 2047;
			 1 : dataOut   <= 2072;
			 2 : dataOut   <= 2097;
			 3 : dataOut   <= 2122;
			 4 : dataOut   <= 2147;
			 5 : dataOut   <= 2173;
			 6 : dataOut   <= 2198;
			 7 : dataOut   <= 2223;
			 8 : dataOut   <= 2248;
			 9 : dataOut   <= 2273;
			10 : dataOut   <= 2298;
			11 : dataOut   <= 2322;
			12 : dataOut   <= 2347;
			13 : dataOut   <= 2372;
			14 : dataOut   <= 2397;
			15 : dataOut   <= 2422;
			16 : dataOut   <= 2446;
			17 : dataOut   <= 2471;
			18 : dataOut   <= 2496;
			19 : dataOut   <= 2520;
			20 : dataOut   <= 2544;
			21 : dataOut   <= 2569;
			22 : dataOut   <= 2593;
			23 : dataOut   <= 2617;
			24 : dataOut   <= 2641;
			25 : dataOut   <= 2665;
			26 : dataOut   <= 2689;
			27 : dataOut   <= 2713;
			28 : dataOut   <= 2737;
			29 : dataOut   <= 2760;
			30 : dataOut   <= 2784;
			31 : dataOut   <= 2807;
			32 : dataOut   <= 2830;
			33 : dataOut   <= 2854;
			34 : dataOut   <= 2877;
			35 : dataOut   <= 2899;
			36 : dataOut   <= 2922;
			37 : dataOut   <= 2945;
			38 : dataOut   <= 2967;
			39 : dataOut   <= 2990;
			40 : dataOut   <= 3012;
			41 : dataOut   <= 3034;
			42 : dataOut   <= 3056;
			43 : dataOut   <= 3078;
			44 : dataOut   <= 3099;
			45 : dataOut   <= 3121;
			46 : dataOut   <= 3142;
			47 : dataOut   <= 3163;
			48 : dataOut   <= 3184;
			49 : dataOut   <= 3205;
			50 : dataOut   <= 3226;
			51 : dataOut   <= 3246;
			52 : dataOut   <= 3266;
			53 : dataOut   <= 3286;
			54 : dataOut   <= 3306;
			55 : dataOut   <= 3326;
			56 : dataOut   <= 3346;
			57 : dataOut   <= 3365;
			58 : dataOut   <= 3384;
			59 : dataOut   <= 3403;
			60 : dataOut   <= 3422;
			61 : dataOut   <= 3440;
			62 : dataOut   <= 3458;
			63 : dataOut   <= 3477;
			64 : dataOut   <= 3494;
			65 : dataOut   <= 3512;
			66 : dataOut   <= 3530;  
			67 : dataOut   <= 3547;
			68 : dataOut   <= 3564;
			69 : dataOut   <= 3580;
			70 : dataOut   <= 3597;
			71 : dataOut   <= 3613;
			72 : dataOut   <= 3629;
			73 : dataOut   <= 3645;
			74 : dataOut   <= 3661;
			75 : dataOut   <= 3676;
			76 : dataOut   <= 3691;
			77 : dataOut   <= 3706;
			78 : dataOut   <= 3721;
			79 : dataOut   <= 3735;
			80 : dataOut   <= 3749;
			81 : dataOut   <= 3763;
			82 : dataOut   <= 3776;
			83 : dataOut   <= 3790;
			84 : dataOut   <= 3803;
			85 : dataOut   <= 3816;
			86 : dataOut   <= 3828;
			87 : dataOut   <= 3840;
			88 : dataOut   <= 3852;
			89 : dataOut   <= 3864;
			90 : dataOut   <= 3875;
			91 : dataOut   <= 3887;
			92 : dataOut   <= 3897;
			93 : dataOut   <= 3908;
			94 : dataOut   <= 3918;
			95 : dataOut   <= 3928;
			96 : dataOut   <= 3938;
			97 : dataOut   <= 3948;
			98 : dataOut   <= 3957;
			99 : dataOut   <= 3966;
			100 : dataOut   <= 3974;
			101 : dataOut   <= 3983;
			102 : dataOut   <= 3991;
			103 : dataOut   <= 3998;
			104 : dataOut   <= 4006;
			105 : dataOut   <= 4013;
			106 : dataOut   <= 4020;
			107 : dataOut   <= 4026;
			108 : dataOut   <= 4033;
			109 : dataOut   <= 4039;
			110 : dataOut   <= 4044;
			111 : dataOut   <= 4050;
			112 : dataOut   <= 4055;
			113 : dataOut   <= 4059;
			114 : dataOut   <= 4064;
			115 : dataOut   <= 4068;
			116 : dataOut   <= 4072;
			117 : dataOut   <= 4075;
			118 : dataOut   <= 4079;
			119 : dataOut   <= 4082;
			120 : dataOut   <= 4084;
			121 : dataOut   <= 4086;
			122 : dataOut   <= 4088;
			123 : dataOut   <= 4090;
			124 : dataOut   <= 4092;
			125 : dataOut   <= 4093;
			126 : dataOut   <= 4093;
			127 : dataOut   <= 4094;
			128 : dataOut   <= 4094;
			129 : dataOut   <= 4094;
			130 : dataOut   <= 4093;
			131 : dataOut   <= 4093;
			132 : dataOut   <= 4092;
			133 : dataOut   <= 4090;
			134 : dataOut   <= 4088;
			135 : dataOut   <= 4086;
			136 : dataOut   <= 4084;
			137 : dataOut   <= 4082;
			138 : dataOut   <= 4079;
			139 : dataOut   <= 4075;
			140 : dataOut   <= 4072;
			141 : dataOut   <= 4068;
			142 : dataOut   <= 4064;
			143 : dataOut   <= 4059;
			144 : dataOut   <= 4055;
			145 : dataOut   <= 4050;
			146 : dataOut   <= 4044;
			147 : dataOut   <= 4039;
			148 : dataOut   <= 4033;
			149 : dataOut   <= 4026;
			150 : dataOut   <= 4020;
			151 : dataOut   <= 4013;
			152 : dataOut   <= 4006;
			153 : dataOut   <= 3998;
			154 : dataOut   <= 3991;
			155 : dataOut   <= 3983;
			156 : dataOut   <= 3974;
			157 : dataOut   <= 3966;
			158 : dataOut   <= 3957;
			159 : dataOut   <= 3948;
			160 : dataOut   <= 3938;
			161 : dataOut   <= 3928;
			162 : dataOut   <= 3918;
			163 : dataOut   <= 3908;
			164 : dataOut   <= 3897;
			165 : dataOut   <= 3887;
			166 : dataOut   <= 3875;
			167 : dataOut   <= 3864;
			168 : dataOut   <= 3852;
			169 : dataOut   <= 3840;
			170 : dataOut   <= 3828;
			171 : dataOut   <= 3816;
			172 : dataOut   <= 3803;
			173 : dataOut   <= 3790;
			174 : dataOut   <= 3776;
			175 : dataOut   <= 3763;
			176 : dataOut   <= 3749;
			177 : dataOut   <= 3735;
			178 : dataOut   <= 3721;
			179 : dataOut   <= 3706;
			180 : dataOut   <= 3691;
			181 : dataOut   <= 3676;
			182 : dataOut   <= 3661;
			183 : dataOut   <= 3645;
			184 : dataOut   <= 3629;
			185 : dataOut   <= 3613;
			186 : dataOut   <= 3597;
			187 : dataOut   <= 3580;
			188 : dataOut   <= 3564;
			189 : dataOut   <= 3547;
			190 : dataOut   <= 3530;
			191 : dataOut   <= 3512;
			192 : dataOut   <= 3494;
			193 : dataOut   <= 3477;
			194 : dataOut   <= 3458;
			195 : dataOut   <= 3440;
			196 : dataOut   <= 3422;
			197 : dataOut   <= 3403;
			198 : dataOut   <= 3384;
			199 : dataOut   <= 3365;
			200 : dataOut   <= 3346;
			201 : dataOut   <= 3326;
			202 : dataOut   <= 3306;
			203 : dataOut   <= 3286;
			204 : dataOut   <= 3266;
			205 : dataOut   <= 3246;
			206 : dataOut   <= 3226;
			207 : dataOut   <= 3205;
			208 : dataOut   <= 3184;
			209 : dataOut   <= 3163;
			210 : dataOut   <= 3142;
			211 : dataOut   <= 3121;
			212 : dataOut   <= 3099;
			213 : dataOut   <= 3078;
			214 : dataOut   <= 3056;
			215 : dataOut   <= 3034;
			216 : dataOut   <= 3012;
			217 : dataOut   <= 2990;
			218 : dataOut   <= 2967;
			219 : dataOut   <= 2945;
			220 : dataOut   <= 2922;
			221 : dataOut   <= 2899;
			222 : dataOut   <= 2877;
			223 : dataOut   <= 2854;
			224 : dataOut   <= 2830;
			225 : dataOut   <= 2807;
			226 : dataOut   <= 2784;
			227 : dataOut   <= 2760;
			228 : dataOut   <= 2737;
			229 : dataOut   <= 2713;
			230 : dataOut   <= 2689;
			231 : dataOut   <= 2665;
			232 : dataOut   <= 2641;
			233 : dataOut   <= 2617;
			234 : dataOut   <= 2593;
			235 : dataOut   <= 2569;
			236 : dataOut   <= 2544;
			237 : dataOut   <= 2520;
			238 : dataOut   <= 2496;
			239 : dataOut   <= 2471;
			240 : dataOut   <= 2446;
			241 : dataOut   <= 2422;
			242 : dataOut   <= 2397;
			243 : dataOut   <= 2372;
			244 : dataOut   <= 2347;
			245 : dataOut   <= 2322;
			246 : dataOut   <= 2298;
			247 : dataOut   <= 2273;
			248 : dataOut   <= 2248;
			249 : dataOut   <= 2223;
			250 : dataOut   <= 2198;
			251 : dataOut   <= 2173;
			252 : dataOut   <= 2147;
			253 : dataOut   <= 2122;
			254 : dataOut   <= 2097;
			255 : dataOut   <= 2072;
			256 : dataOut   <= 2047;
			257 : dataOut   <= 2022;
			258 : dataOut   <= 1997;
			259 : dataOut   <= 1972;
			260 : dataOut   <= 1947;
			261 : dataOut   <= 1921;
			262 : dataOut   <= 1896;
			263 : dataOut   <= 1871;
			264 : dataOut   <= 1846;
			265 : dataOut   <= 1821;
			266 : dataOut   <= 1796;
			267 : dataOut   <= 1772;
			268 : dataOut   <= 1747;
			269 : dataOut   <= 1722;
			270 : dataOut   <= 1697;
			271 : dataOut   <= 1672;
			272 : dataOut   <= 1648;
			273 : dataOut   <= 1623;
			274 : dataOut   <= 1598;
			275 : dataOut   <= 1574;
			276 : dataOut   <= 1550;
			277 : dataOut   <= 1525;
			278 : dataOut   <= 1501;
			279 : dataOut   <= 1477;
			280 : dataOut   <= 1453;
			281 : dataOut   <= 1429;
			282 : dataOut   <= 1405;
			283 : dataOut   <= 1381;
			284 : dataOut   <= 1357;
			285 : dataOut   <= 1334;
			286 : dataOut   <= 1310;
			287 : dataOut   <= 1287;
			288 : dataOut   <= 1264;
			289 : dataOut   <= 1240;
			290 : dataOut   <= 1217;
			291 : dataOut   <= 1195;
			292 : dataOut   <= 1172;
			293 : dataOut   <= 1149;
			294 : dataOut   <= 1127;
			295 : dataOut   <= 1104;
			296 : dataOut   <= 1082;
			297 : dataOut   <= 1060;
			298 : dataOut   <= 1038;
			299 : dataOut   <= 1016;
			300 : dataOut   <= 995;
			301 : dataOut   <= 973;
			302 : dataOut   <= 952;
			303 : dataOut   <= 931;
			304 : dataOut   <= 910;
			305 : dataOut   <= 889;
			306 : dataOut   <= 868;
			307 : dataOut   <= 848;
			308 : dataOut   <= 828;
			309 : dataOut   <= 808;
			310 : dataOut   <= 788;
			311 : dataOut   <= 768;
			312 : dataOut   <= 748;
			313 : dataOut   <= 729;
			314 : dataOut   <= 710;
			315 : dataOut   <= 691;
			316 : dataOut   <= 672;
			317 : dataOut   <= 654;
			318 : dataOut   <= 636;
			319 : dataOut   <= 617;
			320 : dataOut   <= 600;
			321 : dataOut   <= 582;
			322 : dataOut   <= 564;
			323 : dataOut   <= 547;
			324 : dataOut   <= 530;
			325 : dataOut   <= 514;
			326 : dataOut   <= 497;
			327 : dataOut   <= 481;
			328 : dataOut   <= 465;
			329 : dataOut   <= 449;
			330 : dataOut   <= 433;
			331 : dataOut   <= 418;
			332 : dataOut   <= 403;
			333 : dataOut   <= 388;
			334 : dataOut   <= 373;
			335 : dataOut   <= 359;
			336 : dataOut   <= 345;
			337 : dataOut   <= 331;
			338 : dataOut   <= 318;
			339 : dataOut   <= 304;
			340 : dataOut   <= 291;
			341 : dataOut   <= 278;
			342 : dataOut   <= 266;
			343 : dataOut   <= 254;
			344 : dataOut   <= 242;
			345 : dataOut   <= 230;
			346 : dataOut   <= 219;
			347 : dataOut   <= 207;
			348 : dataOut   <= 197;
			349 : dataOut   <= 186;
			350 : dataOut   <= 176;
			351 : dataOut   <= 166;
			352 : dataOut   <= 156;
			353 : dataOut   <= 146;
			354 : dataOut   <= 137;
			355 : dataOut   <= 128;
			356 : dataOut   <= 120;
			357 : dataOut   <= 111;
			358 : dataOut   <= 103;
			359 : dataOut   <= 96;
			360 : dataOut   <= 88;
			361 : dataOut   <= 81;
			362 : dataOut   <= 74;
			363 : dataOut   <= 68;
			364 : dataOut   <= 61;
			365 : dataOut   <= 55;
			366 : dataOut   <= 50;
			367 : dataOut   <= 44;
			368 : dataOut   <= 39;
			369 : dataOut   <= 35;
			370 : dataOut   <= 30;
			371 : dataOut   <= 26;
			372 : dataOut   <= 22;
			373 : dataOut   <= 19;
			374 : dataOut   <= 15;
			375 : dataOut   <= 12;
			376 : dataOut   <= 10;
			377 : dataOut   <= 8;
			378 : dataOut   <= 6;
			379 : dataOut   <= 4;
			380 : dataOut   <= 2;
			381 : dataOut   <= 1;
			382 : dataOut   <= 1;
			383 : dataOut   <= 0;
			384 : dataOut   <= 0;
			385 : dataOut   <= 0;
			386 : dataOut   <= 1;
			387 : dataOut   <= 1;
			388 : dataOut   <= 2;
			389 : dataOut   <= 4;
			390 : dataOut   <= 6;
			391 : dataOut   <= 8;
			392 : dataOut   <= 10;
			393 : dataOut   <= 12;
			394 : dataOut   <= 15;
			395 : dataOut   <= 19;
			396 : dataOut   <= 22;
			397 : dataOut   <= 26;
			398 : dataOut   <= 30;
			399 : dataOut   <= 35;
			400 : dataOut   <= 39;
			401 : dataOut   <= 44;
			402 : dataOut   <= 50;
			403 : dataOut   <= 55;
			404 : dataOut   <= 61;
			405 : dataOut   <= 68;
			406 : dataOut   <= 74;
			407 : dataOut   <= 81;
			408 : dataOut   <= 88;
			409 : dataOut   <= 96;
			410 : dataOut   <= 103;
			411 : dataOut   <= 111;
			412 : dataOut   <= 120;
			413 : dataOut   <= 128;
			414 : dataOut   <= 137;
			415 : dataOut   <= 146;
			416 : dataOut   <= 156;
			417 : dataOut   <= 166;
			418 : dataOut   <= 176;
			419 : dataOut   <= 186;
			420 : dataOut   <= 197;
			421 : dataOut   <= 207;
			422 : dataOut   <= 219;
			423 : dataOut   <= 230;
			424 : dataOut   <= 242;
			425 : dataOut   <= 254;
			426 : dataOut   <= 266;
			427 : dataOut   <= 278;
			428 : dataOut   <= 291;
			429 : dataOut   <= 304;
			430 : dataOut   <= 318;
			431 : dataOut   <= 331;
			432 : dataOut   <= 345;
			433 : dataOut   <= 359;
			434 : dataOut   <= 373;
			435 : dataOut   <= 388;
			436 : dataOut   <= 403;
			437 : dataOut   <= 418;
			438 : dataOut   <= 433;
			439 : dataOut   <= 449;
			440 : dataOut   <= 465;
			441 : dataOut   <= 481;
			442 : dataOut   <= 497;
			443 : dataOut   <= 514;
			444 : dataOut   <= 530;
			445 : dataOut   <= 547;
			446 : dataOut   <= 564;
			447 : dataOut   <= 582;
			448 : dataOut   <= 600;
			449 : dataOut   <= 617;
			450 : dataOut   <= 636;
			451 : dataOut   <= 654;
			452 : dataOut   <= 672;
			453 : dataOut   <= 691;
			454 : dataOut   <= 710;
			455 : dataOut   <= 729;
			456 : dataOut   <= 748;
			457 : dataOut   <= 768;
			458 : dataOut   <= 788;
			459 : dataOut   <= 808;
			460 : dataOut   <= 828;
			461 : dataOut   <= 848;
			462 : dataOut   <= 868;
			463 : dataOut   <= 889;
			464 : dataOut   <= 910;
			465 : dataOut   <= 931;
			466 : dataOut   <= 952;
			467 : dataOut   <= 973;
			468 : dataOut   <= 995;
			469 : dataOut   <= 1016;
			470 : dataOut   <= 1038;
			471 : dataOut   <= 1060;
			472 : dataOut   <= 1082;
			473 : dataOut   <= 1104;
			474 : dataOut   <= 1127;
			475 : dataOut   <= 1149;
			476 : dataOut   <= 1172;
			477 : dataOut   <= 1195;
			478 : dataOut   <= 1217;
			479 : dataOut   <= 1240;
			480 : dataOut   <= 1264;
			481 : dataOut   <= 1287;
			482 : dataOut   <= 1310;
			483 : dataOut   <= 1334;
			484 : dataOut   <= 1357;
			485 : dataOut   <= 1381;
			486 : dataOut   <= 1405;
			487 : dataOut   <= 1429;
			488 : dataOut   <= 1453;
			489 : dataOut   <= 1477;
			490 : dataOut   <= 1501;
			491 : dataOut   <= 1525;
			492 : dataOut   <= 1550;
			493 : dataOut   <= 1574;
			494 : dataOut   <= 1598;
			495 : dataOut   <= 1623;
			496 : dataOut   <= 1648;
			497 : dataOut   <= 1672;
			498 : dataOut   <= 1697;
			499 : dataOut   <= 1722;
			500 : dataOut   <= 1747;
			501 : dataOut   <= 1772;
			502 : dataOut   <= 1796;
			503 : dataOut   <= 1821;
			504 : dataOut   <= 1846;
			505 : dataOut   <= 1871;
			506 : dataOut   <= 1896;
			507 : dataOut   <= 1921;
			508 : dataOut   <= 1947;
			509 : dataOut   <= 1972;
			510 : dataOut   <= 1997;
			511 : dataOut   <= 2022;
	    default:
		       dataOut		<= 0;
    endcase  
  end
*/
  
endmodule
